library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity count1s is
port ( clk    : in      std_ulogic;
       rst_n  : in      std_ulogic;
       onesec_o : out     std_ulogic);
end entity;

architecture rtl of count1s is
  
begin

end architecture rtl;
